.OP
Vs v1 GND 5.248421e+00
R1 v1 v2 1.001471e+03
R2 v3 v2 2.007807e+03
R3 v2 v5 3.112697e+03
R4 v5 GND 4.106096e+03
R5 v5 v6 3.026707e+03
R6 GND v4 2.012925e+03
V6 v4 v7 0.000000e+00
R7 v7 v8 1.029052e+03
C v6 v8 1.040860e-06
Gb v6 v3 v2 v5 7.214136e-03
Hd v5 v8 V6 8.014551e+03
.END
